
module vv 
	input bit A 
	input bit B 
	output bit Q




end module